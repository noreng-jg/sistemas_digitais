LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY converte_neg IS
	PORT(entrada: in std_logic_vector(5 downto 0);  -- entrada binaria
	hex1: out std_logic_vector(6 downto 0); -- saida para o display de sete segmentos
	hex2:out std_logic_vector(6 downto 0);
	hex3:out std_logic_vector(6 downto 0));  
End converte_neg;


architecture sub_arc of converte_neg is 

begin

With entrada select
 hex1 <= "1000000" when "000000" , -- 0
"1111001" when "000001" , -- 1
"0100100" when "000010" , -- 2
"0110000" when "000011" , -- 3
"0011001" when "000100" , -- 4
"0010010" when "000101" , -- 5
"0000010" when "000110" , -- 6
"1111000" when "000111" , -- 7
"0000000" when "001000" , -- 8
"0010000" when "001001" , -- 9
"1000000" when "001010" , -- 0
"1111001" when "001011" , -- 1
"0100100" when "001100" , -- 2
"0110000" when "001101" , -- 3
"0011001" when "001110" , -- 4
"0010010" when "001111" , -- 5
"0000010" when "010000" , -- 6
"1111000" when "010001" , -- 7
"0000000" when "010010" , -- 8
"0010000" when "010011" , -- 9
"1000000" when "010100" , -- 0
"1111001" when "010101" , -- 1
"0100100" when "010110" , -- 2
"0110000" when "010111" , -- 3
"0011001" when "011000" , -- 4
"0010010" when "011001" , -- 5
"0000010" when "011010" , -- 6
"1111000" when "011011" , -- 7
"0000000" when "011100" , -- 8
"0010000" when "011101" , -- 9
"1000000" when "011110" , -- 0
"1111001" when "011111" , -- 1
"0100100" when "100000" , -- 2
"0110000" when "100001" , -- 3
"0011001" when "100010" , -- 4
"0010010" when "100011" , -- 5
"0000010" when "100100" , -- 6
"1111000" when "100101" , -- 7
"0000000" when "100110" , -- 8
"0010000" when "100111" , -- 9
"1000000" when "101000" , -- 0
"1111001" when "101001" , -- 1
"0100100" when "101010" , -- 2
"0110000" when "101011" , -- 3
"0011001" when "101100" , -- 4
"0010010" when "101101" , -- 5
"0000010" when "101110" , -- 6
"1111000" when "101111" , -- 7
"0000000" when "110000" , -- 8
"0010000" when "110001" , -- 9
"1000000" when "110010" , -- 0
"1111001" when "110011" , -- 1
"0100100" when "110100" , -- 2
"0110000" when "110101" , -- 3
"0011001" when "110110" , -- 4
"0010010" when "110111" , -- 5
"0000010" when "111000" , -- 6
"1111000" when "111001" , -- 7
"0000000" when "111010" , -- 8
"0010000" when "111011" , -- 9
"1000000" when "111100" , -- 0
"1111001" when "111101" , -- 1
"0100100" when "111110" , -- 2
"0110000" when "111111" ; -- 3


With entrada select
 hex2 <= "0111111" when "000000" , --   -0
"0111111" when "000001" , --   -0
"0111111" when "000010" , --   -0
"0111111" when "000011" , --   -0
"0111111" when "000100" , --   -0
"0111111" when "000101" , --   -0
"0111111" when "000110" , --   -0
"0111111" when "000111" , --   -0
"0111111" when "001000" , --   -0
"0111111" when "001001" , --   -0
"1111001" when "001010" ,-- %   -10
"1111001" when "001011" ,-- %   -10
"1111001" when "001100" ,-- %   -10
"1111001" when "001101" ,-- %   -10
"1111001" when "001110" ,-- %   -10
"1111001" when "001111" ,-- %   -10
"1111001" when "010000" ,-- %   -10
"1111001" when "010001" ,-- %   -10
"1111001" when "010010" ,-- %   -10
"1111001" when "010011" ,-- %   -10
"0100100" when "010100" ,-- %   -20
"0100100" when "010101" ,-- %   -20
"0100100" when "010110" ,-- %   -20
"0100100" when "010111" ,-- %   -20
"0100100" when "011000" ,-- %   -20
"0100100" when "011001" ,-- %   -20
"0100100" when "011010" ,-- %   -20
"0100100" when "011011" ,-- %   -20
"0100100" when "011100" ,-- %   -20
"0100100" when "011101" ,-- %   -20
"0110000" when "011110" ,-- %   -30
"0110000" when "011111" ,-- %   -30
"0110000" when "100000" ,-- %   -30
"0110000" when "100001" ,-- %   -30
"0110000" when "100010" ,-- %   -30
"0110000" when "100011" ,-- %   -30
"0110000" when "100100" ,-- %   -30
"0110000" when "100101" ,-- %   -30
"0110000" when "100110" ,-- %   -30
"0110000" when "100111" ,-- %   -30
"0011001" when "101000" ,-- %   -40
"0011001" when "101001" ,-- %   -40
"0011001" when "101010" ,-- %   -40
"0011001" when "101011" ,-- %   -40
"0011001" when "101100" ,-- %   -40
"0011001" when "101101" ,-- %   -40
"0011001" when "101110" ,-- %   -40
"0011001" when "101111" ,-- %   -40
"0011001" when "110000" ,-- %   -40
"0011001" when "110001" ,-- %   -40
"0010010" when "110010" ,-- %   -50
"0010010" when "110011" ,-- %   -50
"0010010" when "110100" ,-- %   -50
"0010010" when "110101" ,-- %   -50
"0010010" when "110110" ,-- %   -50
"0010010" when "110111" ,-- %   -50
"0010010" when "111000" ,-- %   -50
"0010010" when "111001" ,-- %   -50
"0010010" when "111010" ,-- %   -50
"0010010" when "111011" ,-- %   -50
"0000010" when "111100" ,-- %   -60
"0000010" when "111101" ,-- %   -60
"0000010" when "111110" ,-- %   -60
"0000010" when "111111" ;-- %   -60


With entrada select
 hex3 <= "1000000" when "000000" ,---   0
"1000000" when "000001" ,---   0
"1000000" when "000010" ,---   0
"1000000" when "000011" ,---   0
"1000000" when "000100" ,---   0
"1000000" when "000101" ,---   0
"1000000" when "000110" ,---   0
"1000000" when "000111" ,---   0
"1000000" when "001000" ,---   0
"1000000" when "001001" ,---   0
"0111111" when "001010" ,---  (-)
"0111111" when "001011" ,---  (-)
"0111111" when "001100" ,---  (-)
"0111111" when "001101" ,---  (-)
"0111111" when "001110" ,---  (-)
"0111111" when "001111" ,---  (-)
"0111111" when "010000" ,---  (-)
"0111111" when "010001" ,---  (-)
"0111111" when "010010" ,---  (-)
"0111111" when "010011" ,---  (-)
"0111111" when "010100" ,---  (-)
"0111111" when "010101" ,---  (-)
"0111111" when "010110" ,---  (-)
"0111111" when "010111" ,---  (-)
"0111111" when "011000" ,---  (-)
"0111111" when "011001" ,---  (-)
"0111111" when "011010" ,---  (-)
"0111111" when "011011" ,---  (-)
"0111111" when "011100" ,---  (-)
"0111111" when "011101" ,---  (-)
"0111111" when "011110" ,---  (-)
"0111111" when "011111" ,---  (-)
"0111111" when "100000" ,---  (-)
"0111111" when "100001" ,---  (-)
"0111111" when "100010" ,---  (-)
"0111111" when "100011" ,---  (-)
"0111111" when "100100" ,---  (-)
"0111111" when "100101" ,---  (-)
"0111111" when "100110" ,---  (-)
"0111111" when "100111" ,---  (-)
"0111111" when "101000" ,---  (-)
"0111111" when "101001" ,---  (-)
"0111111" when "101010" ,---  (-)
"0111111" when "101011" ,---  (-)
"0111111" when "101100" ,---  (-)
"0111111" when "101101" ,---  (-)
"0111111" when "101110" ,---  (-)
"0111111" when "101111" ,---  (-)
"0111111" when "110000" ,---  (-)
"0111111" when "110001" ,---  (-)
"0111111" when "110010" ,---  (-)
"0111111" when "110011" ,---  (-)
"0111111" when "110100" ,---  (-)
"0111111" when "110101" ,---  (-)
"0111111" when "110110" ,---  (-)
"0111111" when "110111" ,---  (-)
"0111111" when "111000" ,---  (-)
"0111111" when "111001" ,---  (-)
"0111111" when "111010" ,---  (-)
"0111111" when "111011" ,---  (-)
"0111111" when "111100" ,---  (-)
"0111111" when "111101" ,---  (-)
"0111111" when "111110" ,---  (-)
"0111111" when "111111" ;---  (-)

end sub_arc;