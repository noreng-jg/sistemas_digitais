LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY converte_soma IS
	PORT(entrada: in std_logic_vector(6 downto 0);  -- entrada binaria
	hex1: out std_logic_vector(6 downto 0); -- saida para o display de sete segmentos
	hex2:out std_logic_vector(6 downto 0); 
	hex3:out std_logic_vector(6 downto 0)); 
End converte_soma;

architecture arc_soma of converte_soma is 
begin

With entrada select
 hex1 <= "1000000" when "0000000" , -- 0
"1111001" when "0000001" , -- 1
"0100100" when "0000010" , -- 2
"0110000" when "0000011" , -- 3
"0011001" when "0000100" , -- 4
"0010010" when "0000101" , -- 5
"0000010" when "0000110" , -- 6
"1111000" when "0000111" , -- 7
"0000000" when "0001000" , -- 8
"0010000" when "0001001" , -- 9
"1000000" when "0001010" , -- 0
"1111001" when "0001011" , -- 1
"0100100" when "0001100" , -- 2
"0110000" when "0001101" , -- 3
"0011001" when "0001110" , -- 4
"0010010" when "0001111" , -- 5
"0000010" when "0010000" , -- 6
"1111000" when "0010001" , -- 7
"0000000" when "0010010" , -- 8
"0010000" when "0010011" , -- 9
"1000000" when "0010100" , -- 0
"1111001" when "0010101" , -- 1
"0100100" when "0010110" , -- 2
"0110000" when "0010111" , -- 3
"0011001" when "0011000" , -- 4
"0010010" when "0011001" , -- 5
"0000010" when "0011010" , -- 6
"1111000" when "0011011" , -- 7
"0000000" when "0011100" , -- 8
"0010000" when "0011101" , -- 9
"1000000" when "0011110" , -- 0
"1111001" when "0011111" , -- 1
"0100100" when "0100000" , -- 2
"0110000" when "0100001" , -- 3
"0011001" when "0100010" , -- 4
"0010010" when "0100011" , -- 5
"0000010" when "0100100" , -- 6
"1111000" when "0100101" , -- 7
"0000000" when "0100110" , -- 8
"0010000" when "0100111" , -- 9
"1000000" when "0101000" , -- 0
"1111001" when "0101001" , -- 1
"0100100" when "0101010" , -- 2
"0110000" when "0101011" , -- 3
"0011001" when "0101100" , -- 4
"0010010" when "0101101" , -- 5
"0000010" when "0101110" , -- 6
"1111000" when "0101111" , -- 7
"0000000" when "0110000" , -- 8
"0010000" when "0110001" , -- 9
"1000000" when "0110010" , -- 0
"1111001" when "0110011" , -- 1
"0100100" when "0110100" , -- 2
"0110000" when "0110101" , -- 3
"0011001" when "0110110" , -- 4
"0010010" when "0110111" , -- 5
"0000010" when "0111000" , -- 6
"1111000" when "0111001" , -- 7
"0000000" when "0111010" , -- 8
"0010000" when "0111011" , -- 9
"1000000" when "0111100" , -- 0
"1111001" when "0111101" , -- 1
"0100100" when "0111110" , -- 2
"0110000" when "0111111" , -- 3
"0011001" when "1000000" , -- 4
"0010010" when "1000001" , -- 5
"0000010" when "1000010" , -- 6
"1111000" when "1000011" , -- 7
"0000000" when "1000100" , -- 8
"0010000" when "1000101" , -- 9
"1000000" when "1000110" , -- 0
"1111001" when "1000111" , -- 1
"0100100" when "1001000" , -- 2
"0110000" when "1001001" , -- 3
"0011001" when "1001010" , -- 4
"0010010" when "1001011" , -- 5
"0000010" when "1001100" , -- 6
"1111000" when "1001101" , -- 7
"0000000" when "1001110" , -- 8
"0010000" when "1001111" , -- 9
"1000000" when "1010000" , -- 0
"1111001" when "1010001" , -- 1
"0100100" when "1010010" , -- 2
"0110000" when "1010011" , -- 3
"0011001" when "1010100" , -- 4
"0010010" when "1010101" , -- 5
"0000010" when "1010110" , -- 6
"1111000" when "1010111" , -- 7
"0000000" when "1011000" , -- 8
"0010000" when "1011001" , -- 9
"1000000" when "1011010" , -- 0
"1111001" when "1011011" , -- 1
"0100100" when "1011100" , -- 2
"0110000" when "1011101" , -- 3
"0011001" when "1011110" , -- 4
"0010010" when "1011111" , -- 5
"0000010" when "1100000" , -- 6
"1111000" when "1100001" , -- 7
"0000000" when "1100010" , -- 8
"0010000" when "1100011" , -- 9
"1000000" when "1100100" , -- 0
"1111001" when "1100101" , -- 1
"0100100" when "1100110" , -- 2
"0110000" when "1100111" , -- 3
"0011001" when "1101000" , -- 4
"0010010" when "1101001" , -- 5
"0000010" when "1101010" , -- 6
"1111000" when "1101011" , -- 7
"0000000" when "1101100" , -- 8
"0010000" when "1101101" , -- 9
"1000000" when "1101110" , -- 0
"1111001" when "1101111" , -- 1
"0100100" when "1110000" , -- 2
"0110000" when "1110001" , -- 3
"0011001" when "1110010" , -- 4
"0010010" when "1110011" , -- 5
"0000010" when "1110100" , -- 6
"1111000" when "1110101" , -- 7
"0000000" when "1110110" , -- 8
"0010000" when "1110111" , -- 9
"1000000" when "1111000" , -- 0
"1111001" when "1111001" , -- 1
"0100100" when "1111010" , -- 2
"0110000" when "1111011" , -- 3
"0011001" when "1111100" , -- 4
"0010010" when "1111101" , -- 5
"0000010" when "1111110" , -- 6
"1111000" when "1111111" ; --7


With entrada select
 hex2 <= "1000000" when "0000000" , -- 0
"1000000" when "0000001" , -- 0
"1000000" when "0000010" , -- 0
"1000000" when "0000011" , -- 0
"1000000" when "0000100" , -- 0
"1000000" when "0000101" , -- 0
"1000000" when "0000110" , -- 0
"1000000" when "0000111" , -- 0
"1000000" when "0001000" , -- 0
"1000000" when "0001001" , -- 0
"1111001" when "0001010" , -- 10
"1111001" when "0001011" , -- 10
"1111001" when "0001100" , -- 10
"1111001" when "0001101" , -- 10
"1111001" when "0001110" , -- 10
"1111001" when "0001111" , -- 10
"1111001" when "0010000" , -- 10
"1111001" when "0010001" , -- 10
"1111001" when "0010010" , -- 10
"1111001" when "0010011" , -- 10
"0100100" when "0010100" , -- 20
"0100100" when "0010101" , -- 20
"0100100" when "0010110" , -- 20
"0100100" when "0010111" , -- 20
"0100100" when "0011000" , -- 20
"0100100" when "0011001" , -- 20
"0100100" when "0011010" , -- 20
"0100100" when "0011011" , -- 20
"0100100" when "0011100" , -- 20
"0100100" when "0011101" , -- 20
"0110000" when "0011110" , -- 30
"0110000" when "0011111" , -- 30
"0110000" when "0100000" , -- 30
"0110000" when "0100001" , -- 30
"0110000" when "0100010" , -- 30
"0110000" when "0100011" , -- 30
"0110000" when "0100100" , -- 30
"0110000" when "0100101" , -- 30
"0110000" when "0100110" , -- 30
"0110000" when "0100111" , -- 30
"0011001" when "0101000" , -- 40
"0011001" when "0101001" , -- 40
"0011001" when "0101010" , -- 40
"0011001" when "0101011" , -- 40
"0011001" when "0101100" , -- 40
"0011001" when "0101101" , -- 40
"0011001" when "0101110" , -- 40
"0011001" when "0101111" , -- 40
"0011001" when "0110000" , -- 40
"0011001" when "0110001" , -- 40
"0010010" when "0110010" , -- 50
"0010010" when "0110011" , -- 50
"0010010" when "0110100" , -- 50
"0010010" when "0110101" , -- 50
"0010010" when "0110110" , -- 50
"0010010" when "0110111" , -- 50
"0010010" when "0111000" , -- 50
"0010010" when "0111001" , -- 50
"0010010" when "0111010" , -- 50
"0010010" when "0111011" , -- 50
"0000010" when "0111100" , -- 60
"0000010" when "0111101" , -- 60
"0000010" when "0111110" , -- 60
"0000010" when "0111111" , -- 60
"0000010" when "1000000" , -- 60
"0000010" when "1000001" , -- 60
"0000010" when "1000010" , -- 60
"0000010" when "1000011" , -- 60
"0000010" when "1000100" , -- 60
"0000010" when "1000101" , -- 60
"1111000" when "1000110" , -- 70
"1111000" when "1000111" , -- 70
"1111000" when "1001000" , -- 70
"1111000" when "1001001" , -- 70
"1111000" when "1001010" , -- 70
"1111000" when "1001011" , -- 70
"1111000" when "1001100" , -- 70
"1111000" when "1001101" , -- 70
"1111000" when "1001110" , -- 70
"1111000" when "1001111" , -- 70
"0000000" when "1010000" , -- 80
"0000000" when "1010001" , -- 80
"0000000" when "1010010" , -- 80
"0000000" when "1010011" , -- 80
"0000000" when "1010100" , -- 80
"0000000" when "1010101" , -- 80
"0000000" when "1010110" , -- 80
"0000000" when "1010111" , -- 80
"0000000" when "1011000" , -- 80
"0000000" when "1011001" , -- 80
"0010000" when "1011010" , -- 90
"0010000" when "1011011" , -- 90
"0010000" when "1011100" , -- 90
"0010000" when "1011101" , -- 90
"0010000" when "1011110" , -- 90
"0010000" when "1011111" , -- 90
"0010000" when "1100000" , -- 90
"0010000" when "1100001" , -- 90
"0010000" when "1100010" , -- 90
"0010000" when "1100011" , -- 90
"1000000" when "1100100" , -- 0
"1000000" when "1100101" , -- 0
"1000000" when "1100110" , -- 0
"1000000" when "1100111" , -- 0
"1000000" when "1101000" , -- 0
"1000000" when "1101001" , -- 0
"1000000" when "1101010" , -- 0
"1000000" when "1101011" , -- 0
"1000000" when "1101100" , -- 0
"1000000" when "1101101" , -- 0
"1111001" when "1101110" , -- 10
"1111001" when "1101111" , -- 10
"1111001" when "1110000" , -- 10
"1111001" when "1110001" , -- 10
"1111001" when "1110010" , -- 10
"1111001" when "1110011" , -- 10
"1111001" when "1110100" , -- 10
"1111001" when "1110101" , -- 10
"1111001" when "1110110" , -- 10
"1111001" when "1110111" , -- 10
"0100100" when "1111000" , -- 20
"0100100" when "1111001" , -- 20
"0100100" when "1111010" , -- 20
"0100100" when "1111011" , -- 20
"0100100" when "1111100" , -- 20
"0100100" when "1111101" , -- 20
"0100100" when "1111110" , -- 20
"0100100" when "1111111" ; -- 20


With entrada select
 hex3 <= "1000000" when "0000000" , --0 
"1000000" when "0000001" , --0 
"1000000" when "0000010" , --0 
"1000000" when "0000011" , --0 
"1000000" when "0000100" , --0 
"1000000" when "0000101" , --0 
"1000000" when "0000110" , --0 
"1000000" when "0000111" , --0 
"1000000" when "0001000" , --0 
"1000000" when "0001001" , --0 
"1000000" when "0001010" , --0 
"1000000" when "0001011" , --0 
"1000000" when "0001100" , --0 
"1000000" when "0001101" , --0 
"1000000" when "0001110" , --0 
"1000000" when "0001111" , --0 
"1000000" when "0010000" , --0 
"1000000" when "0010001" , --0 
"1000000" when "0010010" , --0 
"1000000" when "0010011" , --0 
"1000000" when "0010100" , --0 
"1000000" when "0010101" , --0 
"1000000" when "0010110" , --0 
"1000000" when "0010111" , --0 
"1000000" when "0011000" , --0 
"1000000" when "0011001" , --0 
"1000000" when "0011010" , --0 
"1000000" when "0011011" , --0 
"1000000" when "0011100" , --0 
"1000000" when "0011101" , --0 
"1000000" when "0011110" , --0 
"1000000" when "0011111" , --0 
"1000000" when "0100000" , --0 
"1000000" when "0100001" , --0 
"1000000" when "0100010" , --0 
"1000000" when "0100011" , --0 
"1000000" when "0100100" , --0 
"1000000" when "0100101" , --0 
"1000000" when "0100110" , --0 
"1000000" when "0100111" , --0 
"1000000" when "0101000" , --0 
"1000000" when "0101001" , --0 
"1000000" when "0101010" , --0 
"1000000" when "0101011" , --0 
"1000000" when "0101100" , --0 
"1000000" when "0101101" , --0 
"1000000" when "0101110" , --0 
"1000000" when "0101111" , --0 
"1000000" when "0110000" , --0 
"1000000" when "0110001" , --0 
"1000000" when "0110010" , --0 
"1000000" when "0110011" , --0 
"1000000" when "0110100" , --0 
"1000000" when "0110101" , --0 
"1000000" when "0110110" , --0 
"1000000" when "0110111" , --0 
"1000000" when "0111000" , --0 
"1000000" when "0111001" , --0 
"1000000" when "0111010" , --0 
"1000000" when "0111011" , --0 
"1000000" when "0111100" , --0 
"1000000" when "0111101" , --0 
"1000000" when "0111110" , --0 
"1000000" when "0111111" , --0 
"1000000" when "1000000" , --0 
"1000000" when "1000001" , --0 
"1000000" when "1000010" , --0 
"1000000" when "1000011" , --0 
"1000000" when "1000100" , --0 
"1000000" when "1000101" , --0 
"1000000" when "1000110" , --0 
"1000000" when "1000111" , --0 
"1000000" when "1001000" , --0 
"1000000" when "1001001" , --0 
"1000000" when "1001010" , --0 
"1000000" when "1001011" , --0 
"1000000" when "1001100" , --0 
"1000000" when "1001101" , --0 
"1000000" when "1001110" , --0 
"1000000" when "1001111" , --0 
"1000000" when "1010000" , --0 
"1000000" when "1010001" , --0 
"1000000" when "1010010" , --0 
"1000000" when "1010011" , --0 
"1000000" when "1010100" , --0 
"1000000" when "1010101" , --0 
"1000000" when "1010110" , --0 
"1000000" when "1010111" , --0 
"1000000" when "1011000" , --0 
"1000000" when "1011001" , --0 
"1000000" when "1011010" , --0 
"1000000" when "1011011" , --0 
"1000000" when "1011100" , --0 
"1000000" when "1011101" , --0 
"1000000" when "1011110" , --0 
"1000000" when "1011111" , --0 
"1000000" when "1100000" , --0 
"1000000" when "1100001" , --0 
"1000000" when "1100010" , --0 
"1000000" when "1100011" , --0 
"1111001" when "1100100" , --100 
"1111001" when "1100101" , --100 
"1111001" when "1100110" , --100 
"1111001" when "1100111" , --100 
"1111001" when "1101000" , --100 
"1111001" when "1101001" , --100 
"1111001" when "1101010" , --100 
"1111001" when "1101011" , --100 
"1111001" when "1101100" , --100 
"1111001" when "1101101" , --100 
"1111001" when "1101110" , --100 
"1111001" when "1101111" , --100 
"1111001" when "1110000" , --100 
"1111001" when "1110001" , --100 
"1111001" when "1110010" , --100 
"1111001" when "1110011" , --100 
"1111001" when "1110100" , --100 
"1111001" when "1110101" , --100 
"1111001" when "1110110" , --100 
"1111001" when "1110111" , --100 
"1111001" when "1111000" , --100 
"1111001" when "1111001" , --100 
"1111001" when "1111010" , --100 
"1111001" when "1111011" , --100 
"1111001" when "1111100" , --100 
"1111001" when "1111101" , --100 
"1111001" when "1111110" , --100 
"1111001" when "1111111" ; --100

end arc_soma;